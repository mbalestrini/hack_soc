VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRF_2R1W
  CLASS BLOCK ;
  FOREIGN DFFRF_2R1W ;
  ORIGIN 0.000 0.000 ;
  SIZE 378.700 BY 176.800 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.830 2.450 ;
    END
  END CLK
  PIN DA[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 0.000 0.690 10.240 ;
    END
  END DA[0]
  PIN DA[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.510 6.020 ;
    END
  END DA[10]
  PIN DA[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.030 2.280 ;
    END
  END DA[11]
  PIN DA[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.090 3.130 ;
    END
  END DA[12]
  PIN DA[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.610 3.130 ;
    END
  END DA[13]
  PIN DA[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.130 9.900 ;
    END
  END DA[14]
  PIN DA[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.190 9.900 ;
    END
  END DA[15]
  PIN DA[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.710 7.180 ;
    END
  END DA[16]
  PIN DA[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.230 2.920 ;
    END
  END DA[17]
  PIN DA[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.750 3.810 ;
    END
  END DA[18]
  PIN DA[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.810 2.280 ;
    END
  END DA[19]
  PIN DA[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.750 8.360 ;
    END
  END DA[1]
  PIN DA[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.330 20.810 ;
    END
  END DA[20]
  PIN DA[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.850 24.210 ;
    END
  END DA[21]
  PIN DA[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.370 2.450 ;
    END
  END DA[22]
  PIN DA[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.430 2.280 ;
    END
  END DA[23]
  PIN DA[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 129.950 5.850 ;
    END
  END DA[24]
  PIN DA[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.470 9.720 ;
    END
  END DA[25]
  PIN DA[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 140.990 7.210 ;
    END
  END DA[26]
  PIN DA[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.050 14.010 ;
    END
  END DA[27]
  PIN DA[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.570 2.280 ;
    END
  END DA[28]
  PIN DA[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.090 3.130 ;
    END
  END DA[29]
  PIN DA[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.270 16.050 ;
    END
  END DA[2]
  PIN DA[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.150 5.170 ;
    END
  END DA[30]
  PIN DA[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.670 24.040 ;
    END
  END DA[31]
  PIN DA[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.790 34.240 ;
    END
  END DA[3]
  PIN DA[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.850 3.300 ;
    END
  END DA[4]
  PIN DA[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.370 20.600 ;
    END
  END DA[5]
  PIN DA[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 32.890 23.530 ;
    END
  END DA[6]
  PIN DA[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.410 4.800 ;
    END
  END DA[7]
  PIN DA[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.470 18.260 ;
    END
  END DA[8]
  PIN DA[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 48.990 15.680 ;
    END
  END DA[9]
  PIN DB[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 173.020 2.530 176.800 ;
    END
  END DB[0]
  PIN DB[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 174.350 93.610 176.800 ;
    END
  END DB[10]
  PIN DB[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 54.020 102.810 176.800 ;
    END
  END DB[11]
  PIN DB[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 172.820 112.010 176.800 ;
    END
  END DB[12]
  PIN DB[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 174.520 120.750 176.800 ;
    END
  END DB[13]
  PIN DB[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 174.520 129.950 176.800 ;
    END
  END DB[14]
  PIN DB[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 170.270 139.150 176.800 ;
    END
  END DB[15]
  PIN DB[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 174.520 148.350 176.800 ;
    END
  END DB[16]
  PIN DB[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 174.520 157.550 176.800 ;
    END
  END DB[17]
  PIN DB[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 174.350 166.750 176.800 ;
    END
  END DB[18]
  PIN DB[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 174.520 175.490 176.800 ;
    END
  END DB[19]
  PIN DB[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 173.360 11.270 176.800 ;
    END
  END DB[1]
  PIN DB[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 158.400 184.690 176.800 ;
    END
  END DB[20]
  PIN DB[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 160.100 193.890 176.800 ;
    END
  END DB[21]
  PIN DB[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 174.520 203.090 176.800 ;
    END
  END DB[22]
  PIN DB[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 174.520 212.290 176.800 ;
    END
  END DB[23]
  PIN DB[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 174.520 221.490 176.800 ;
    END
  END DB[24]
  PIN DB[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 174.520 230.230 176.800 ;
    END
  END DB[25]
  PIN DB[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 174.520 239.430 176.800 ;
    END
  END DB[26]
  PIN DB[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 174.520 248.630 176.800 ;
    END
  END DB[27]
  PIN DB[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 165.510 257.830 176.800 ;
    END
  END DB[28]
  PIN DB[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 170.980 267.030 176.800 ;
    END
  END DB[29]
  PIN DB[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 174.350 20.470 176.800 ;
    END
  END DB[2]
  PIN DB[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 173.020 276.230 176.800 ;
    END
  END DB[30]
  PIN DB[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 173.360 284.970 176.800 ;
    END
  END DB[31]
  PIN DB[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 146.500 29.670 176.800 ;
    END
  END DB[3]
  PIN DB[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 163.680 38.870 176.800 ;
    END
  END DB[4]
  PIN DB[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 174.350 48.070 176.800 ;
    END
  END DB[5]
  PIN DB[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 126.280 57.270 176.800 ;
    END
  END DB[6]
  PIN DB[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 174.350 66.010 176.800 ;
    END
  END DB[7]
  PIN DB[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 166.870 75.210 176.800 ;
    END
  END DB[8]
  PIN DB[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 157.380 84.410 176.800 ;
    END
  END DB[9]
  PIN DW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.190 6.320 ;
    END
  END DW[0]
  PIN DW[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 0.000 227.010 4.460 ;
    END
  END DW[10]
  PIN DW[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.530 24.000 ;
    END
  END DW[11]
  PIN DW[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.050 21.960 ;
    END
  END DW[12]
  PIN DW[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.110 25.570 ;
    END
  END DW[13]
  PIN DW[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.630 2.280 ;
    END
  END DW[14]
  PIN DW[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.150 2.280 ;
    END
  END DW[15]
  PIN DW[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.670 3.980 ;
    END
  END DW[16]
  PIN DW[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.730 2.450 ;
    END
  END DW[17]
  PIN DW[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.250 2.450 ;
    END
  END DW[18]
  PIN DW[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.770 28.760 ;
    END
  END DW[19]
  PIN DW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.710 4.320 ;
    END
  END DW[1]
  PIN DW[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.290 42.540 ;
    END
  END DW[20]
  PIN DW[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.350 37.100 ;
    END
  END DW[21]
  PIN DW[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 291.870 2.450 ;
    END
  END DW[22]
  PIN DW[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.390 13.870 ;
    END
  END DW[23]
  PIN DW[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 302.910 15.680 ;
    END
  END DW[24]
  PIN DW[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 307.970 2.450 ;
    END
  END DW[25]
  PIN DW[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.490 2.450 ;
    END
  END DW[26]
  PIN DW[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.010 2.450 ;
    END
  END DW[27]
  PIN DW[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.070 37.440 ;
    END
  END DW[28]
  PIN DW[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.590 21.120 ;
    END
  END DW[29]
  PIN DW[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.770 8.570 ;
    END
  END DW[2]
  PIN DW[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.110 18.400 ;
    END
  END DW[30]
  PIN DW[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.630 13.870 ;
    END
  END DW[31]
  PIN DW[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.290 2.450 ;
    END
  END DW[3]
  PIN DW[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.810 40.320 ;
    END
  END DW[4]
  PIN DW[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.330 10.240 ;
    END
  END DW[5]
  PIN DW[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.390 24.210 ;
    END
  END DW[6]
  PIN DW[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 0.000 210.910 10.240 ;
    END
  END DW[7]
  PIN DW[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.430 32.160 ;
    END
  END DW[8]
  PIN DW[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 221.950 17.410 ;
    END
  END DW[9]
  PIN RA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.690 24.860 ;
    END
  END RA[0]
  PIN RA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.210 5.850 ;
    END
  END RA[1]
  PIN RA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.730 8.880 ;
    END
  END RA[2]
  PIN RA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.250 12.650 ;
    END
  END RA[3]
  PIN RA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.310 14.660 ;
    END
  END RA[4]
  PIN RB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 168.260 294.170 176.800 ;
    END
  END RB[0]
  PIN RB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 153.480 303.370 176.800 ;
    END
  END RB[1]
  PIN RB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 158.400 312.570 176.800 ;
    END
  END RB[2]
  PIN RB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 157.380 321.770 176.800 ;
    END
  END RB[3]
  PIN RB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 80.510 330.970 176.800 ;
    END
  END RB[4]
  PIN RW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 174.560 339.710 176.800 ;
    END
  END RW[0]
  PIN RW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 150.080 348.910 176.800 ;
    END
  END RW[1]
  PIN RW[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 149.020 358.110 176.800 ;
    END
  END RW[2]
  PIN RW[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 156.200 367.310 176.800 ;
    END
  END RW[3]
  PIN RW[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 156.020 376.510 176.800 ;
    END
  END RW[4]
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.850 136.835 378.510 138.435 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.850 36.835 378.510 38.435 ;
    END
  END VPWR
  PIN WE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.350 17.040 ;
    END
  END WE
  OBS
      LAYER li1 ;
        RECT 0.075 0.085 378.510 176.715 ;
      LAYER met1 ;
        RECT 0.000 0.040 378.510 176.760 ;
      LAYER met2 ;
        RECT 0.030 172.740 2.110 176.790 ;
        RECT 2.810 173.080 10.850 176.790 ;
        RECT 11.550 174.070 20.050 176.790 ;
        RECT 20.750 174.070 29.250 176.790 ;
        RECT 11.550 173.080 29.250 174.070 ;
        RECT 2.810 172.740 29.250 173.080 ;
        RECT 0.030 146.220 29.250 172.740 ;
        RECT 29.950 163.400 38.450 176.790 ;
        RECT 39.150 174.070 47.650 176.790 ;
        RECT 48.350 174.070 56.850 176.790 ;
        RECT 39.150 163.400 56.850 174.070 ;
        RECT 29.950 146.220 56.850 163.400 ;
        RECT 0.030 126.000 56.850 146.220 ;
        RECT 57.550 174.070 65.590 176.790 ;
        RECT 66.290 174.070 74.790 176.790 ;
        RECT 57.550 166.590 74.790 174.070 ;
        RECT 75.490 166.590 83.990 176.790 ;
        RECT 57.550 157.100 83.990 166.590 ;
        RECT 84.690 174.070 93.190 176.790 ;
        RECT 93.890 174.070 102.390 176.790 ;
        RECT 84.690 157.100 102.390 174.070 ;
        RECT 57.550 126.000 102.390 157.100 ;
        RECT 0.030 53.740 102.390 126.000 ;
        RECT 103.090 172.540 111.590 176.790 ;
        RECT 112.290 174.240 120.330 176.790 ;
        RECT 121.030 174.240 129.530 176.790 ;
        RECT 130.230 174.240 138.730 176.790 ;
        RECT 112.290 172.540 138.730 174.240 ;
        RECT 103.090 169.990 138.730 172.540 ;
        RECT 139.430 174.240 147.930 176.790 ;
        RECT 148.630 174.240 157.130 176.790 ;
        RECT 157.830 174.240 166.330 176.790 ;
        RECT 139.430 174.070 166.330 174.240 ;
        RECT 167.030 174.240 175.070 176.790 ;
        RECT 175.770 174.240 184.270 176.790 ;
        RECT 167.030 174.070 184.270 174.240 ;
        RECT 139.430 169.990 184.270 174.070 ;
        RECT 103.090 158.120 184.270 169.990 ;
        RECT 184.970 159.820 193.470 176.790 ;
        RECT 194.170 174.240 202.670 176.790 ;
        RECT 203.370 174.240 211.870 176.790 ;
        RECT 212.570 174.240 221.070 176.790 ;
        RECT 221.770 174.240 229.810 176.790 ;
        RECT 230.510 174.240 239.010 176.790 ;
        RECT 239.710 174.240 248.210 176.790 ;
        RECT 248.910 174.240 257.410 176.790 ;
        RECT 194.170 165.230 257.410 174.240 ;
        RECT 258.110 170.700 266.610 176.790 ;
        RECT 267.310 172.740 275.810 176.790 ;
        RECT 276.510 173.080 284.550 176.790 ;
        RECT 285.250 173.080 293.750 176.790 ;
        RECT 276.510 172.740 293.750 173.080 ;
        RECT 267.310 170.700 293.750 172.740 ;
        RECT 258.110 167.980 293.750 170.700 ;
        RECT 294.450 167.980 302.950 176.790 ;
        RECT 258.110 165.230 302.950 167.980 ;
        RECT 194.170 159.820 302.950 165.230 ;
        RECT 184.970 158.120 302.950 159.820 ;
        RECT 103.090 153.200 302.950 158.120 ;
        RECT 303.650 158.120 312.150 176.790 ;
        RECT 312.850 158.120 321.350 176.790 ;
        RECT 303.650 157.100 321.350 158.120 ;
        RECT 322.050 157.100 330.550 176.790 ;
        RECT 303.650 153.200 330.550 157.100 ;
        RECT 103.090 80.230 330.550 153.200 ;
        RECT 331.250 174.280 339.290 176.790 ;
        RECT 339.990 174.280 348.490 176.790 ;
        RECT 331.250 149.800 348.490 174.280 ;
        RECT 349.190 149.800 357.690 176.790 ;
        RECT 331.250 148.740 357.690 149.800 ;
        RECT 358.390 155.920 366.890 176.790 ;
        RECT 367.590 155.920 376.090 176.790 ;
        RECT 358.390 155.740 376.090 155.920 ;
        RECT 376.790 155.740 378.410 176.790 ;
        RECT 358.390 148.740 378.410 155.740 ;
        RECT 331.250 80.230 378.410 148.740 ;
        RECT 103.090 53.740 378.410 80.230 ;
        RECT 0.030 42.820 378.410 53.740 ;
        RECT 0.030 40.600 280.870 42.820 ;
        RECT 0.030 34.520 194.390 40.600 ;
        RECT 0.030 16.330 16.370 34.520 ;
        RECT 0.030 10.520 10.850 16.330 ;
        RECT 0.030 0.010 0.270 10.520 ;
        RECT 0.970 8.640 10.850 10.520 ;
        RECT 0.970 0.010 5.330 8.640 ;
        RECT 6.030 0.010 10.850 8.640 ;
        RECT 11.550 0.010 16.370 16.330 ;
        RECT 17.070 24.490 194.390 34.520 ;
        RECT 17.070 23.810 113.430 24.490 ;
        RECT 17.070 20.880 32.470 23.810 ;
        RECT 17.070 3.580 26.950 20.880 ;
        RECT 17.070 0.010 21.430 3.580 ;
        RECT 22.130 0.010 26.950 3.580 ;
        RECT 27.650 0.010 32.470 20.880 ;
        RECT 33.170 21.090 113.430 23.810 ;
        RECT 33.170 18.540 107.910 21.090 ;
        RECT 33.170 5.080 43.050 18.540 ;
        RECT 33.170 0.010 37.990 5.080 ;
        RECT 38.690 0.010 43.050 5.080 ;
        RECT 43.750 15.960 107.910 18.540 ;
        RECT 43.750 0.010 48.570 15.960 ;
        RECT 49.270 10.180 107.910 15.960 ;
        RECT 49.270 6.300 75.710 10.180 ;
        RECT 49.270 0.010 54.090 6.300 ;
        RECT 54.790 3.410 75.710 6.300 ;
        RECT 54.790 2.560 64.670 3.410 ;
        RECT 54.790 0.010 59.610 2.560 ;
        RECT 60.310 0.010 64.670 2.560 ;
        RECT 65.370 0.010 70.190 3.410 ;
        RECT 70.890 0.010 75.710 3.410 ;
        RECT 76.410 0.010 80.770 10.180 ;
        RECT 81.470 7.460 107.910 10.180 ;
        RECT 81.470 0.010 86.290 7.460 ;
        RECT 86.990 4.090 107.910 7.460 ;
        RECT 86.990 3.200 97.330 4.090 ;
        RECT 86.990 0.010 91.810 3.200 ;
        RECT 92.510 0.010 97.330 3.200 ;
        RECT 98.030 2.560 107.910 4.090 ;
        RECT 98.030 0.010 102.390 2.560 ;
        RECT 103.090 0.010 107.910 2.560 ;
        RECT 108.610 0.010 113.430 21.090 ;
        RECT 114.130 24.320 194.390 24.490 ;
        RECT 114.130 14.290 167.250 24.320 ;
        RECT 114.130 10.000 145.630 14.290 ;
        RECT 114.130 6.130 135.050 10.000 ;
        RECT 114.130 2.730 129.530 6.130 ;
        RECT 114.130 0.010 118.950 2.730 ;
        RECT 119.650 2.560 129.530 2.730 ;
        RECT 119.650 0.010 124.010 2.560 ;
        RECT 124.710 0.010 129.530 2.560 ;
        RECT 130.230 0.010 135.050 6.130 ;
        RECT 135.750 7.490 145.630 10.000 ;
        RECT 135.750 0.010 140.570 7.490 ;
        RECT 141.270 0.010 145.630 7.490 ;
        RECT 146.330 5.450 167.250 14.290 ;
        RECT 146.330 3.410 161.730 5.450 ;
        RECT 146.330 2.560 156.670 3.410 ;
        RECT 146.330 0.010 151.150 2.560 ;
        RECT 151.850 0.010 156.670 2.560 ;
        RECT 157.370 0.010 161.730 3.410 ;
        RECT 162.430 0.010 167.250 5.450 ;
        RECT 167.950 8.850 194.390 24.320 ;
        RECT 167.950 6.600 183.350 8.850 ;
        RECT 167.950 0.010 172.770 6.600 ;
        RECT 173.470 4.600 183.350 6.600 ;
        RECT 173.470 0.010 178.290 4.600 ;
        RECT 178.990 0.010 183.350 4.600 ;
        RECT 184.050 2.730 194.390 8.850 ;
        RECT 184.050 0.010 188.870 2.730 ;
        RECT 189.570 0.010 194.390 2.730 ;
        RECT 195.090 32.440 280.870 40.600 ;
        RECT 195.090 24.490 216.010 32.440 ;
        RECT 195.090 10.520 204.970 24.490 ;
        RECT 195.090 0.010 199.910 10.520 ;
        RECT 200.610 0.010 204.970 10.520 ;
        RECT 205.670 10.520 216.010 24.490 ;
        RECT 205.670 0.010 210.490 10.520 ;
        RECT 211.190 0.010 216.010 10.520 ;
        RECT 216.710 29.040 280.870 32.440 ;
        RECT 216.710 25.850 275.350 29.040 ;
        RECT 216.710 24.280 242.690 25.850 ;
        RECT 216.710 17.690 232.110 24.280 ;
        RECT 216.710 0.010 221.530 17.690 ;
        RECT 222.230 4.740 232.110 17.690 ;
        RECT 222.230 0.010 226.590 4.740 ;
        RECT 227.290 0.010 232.110 4.740 ;
        RECT 232.810 22.240 242.690 24.280 ;
        RECT 232.810 0.010 237.630 22.240 ;
        RECT 238.330 0.010 242.690 22.240 ;
        RECT 243.390 4.260 275.350 25.850 ;
        RECT 243.390 2.560 259.250 4.260 ;
        RECT 243.390 0.010 248.210 2.560 ;
        RECT 248.910 0.010 253.730 2.560 ;
        RECT 254.430 0.010 259.250 2.560 ;
        RECT 259.950 2.730 275.350 4.260 ;
        RECT 259.950 0.010 264.310 2.730 ;
        RECT 265.010 0.010 269.830 2.730 ;
        RECT 270.530 0.010 275.350 2.730 ;
        RECT 276.050 0.010 280.870 29.040 ;
        RECT 281.570 37.720 378.410 42.820 ;
        RECT 281.570 37.380 323.650 37.720 ;
        RECT 281.570 0.010 285.930 37.380 ;
        RECT 286.630 15.960 323.650 37.380 ;
        RECT 286.630 14.150 302.490 15.960 ;
        RECT 286.630 2.730 296.970 14.150 ;
        RECT 286.630 0.010 291.450 2.730 ;
        RECT 292.150 0.010 296.970 2.730 ;
        RECT 297.670 0.010 302.490 14.150 ;
        RECT 303.190 2.730 323.650 15.960 ;
        RECT 303.190 0.010 307.550 2.730 ;
        RECT 308.250 0.010 313.070 2.730 ;
        RECT 313.770 0.010 318.590 2.730 ;
        RECT 319.290 0.010 323.650 2.730 ;
        RECT 324.350 25.140 378.410 37.720 ;
        RECT 324.350 21.400 345.270 25.140 ;
        RECT 324.350 0.010 329.170 21.400 ;
        RECT 329.870 18.680 345.270 21.400 ;
        RECT 329.870 0.010 334.690 18.680 ;
        RECT 335.390 14.150 345.270 18.680 ;
        RECT 335.390 0.010 340.210 14.150 ;
        RECT 340.910 0.010 345.270 14.150 ;
        RECT 345.970 17.320 378.410 25.140 ;
        RECT 345.970 14.940 377.930 17.320 ;
        RECT 345.970 12.930 366.890 14.940 ;
        RECT 345.970 9.160 361.830 12.930 ;
        RECT 345.970 6.130 356.310 9.160 ;
        RECT 345.970 0.010 350.790 6.130 ;
        RECT 351.490 0.010 356.310 6.130 ;
        RECT 357.010 0.010 361.830 9.160 ;
        RECT 362.530 0.010 366.890 12.930 ;
        RECT 367.590 2.730 377.930 14.940 ;
        RECT 367.590 0.010 372.410 2.730 ;
        RECT 373.110 0.010 377.930 2.730 ;
      LAYER met3 ;
        RECT 1.835 138.835 376.605 176.625 ;
        RECT 1.835 38.835 376.605 136.435 ;
        RECT 1.835 0.175 376.605 36.435 ;
  END
END DFFRF_2R1W
END LIBRARY

