`default_nettype none
`timescale 1ns/10ps

module device_mgr(
	
);

endmodule